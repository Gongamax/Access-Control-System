library ieee;
use ieee.std_logic_1164.all;

entity RingBufferControl is 
Port(--Input ports
     DAV		: in std_logic;
     CTS			: in std_logic;
	  full		: in std_logic;
	  empty		: in std_logic;
	  clk			: in std_logic;
	  reset		: in std_logic;
	  --Output ports
	  Wr		   : out std_logic;
	  selnPG		: out std_logic;
	  incPut		: out std_logic;
	  incGet		: out std_logic;
	  Wreg		: out std_logic;
	  DAC			: out std_logic
);
	  
end RingBufferControl;

architecture behavioral of RingBufferControl is

type State is (Start, Write_memory, Write_done, IncrPut, Finish_write, Attend_output, Output_done);

signal CurrentState, NextState : State;

begin
CurrentState <= Start when reset = '1' else NextState when rising_edge(clk);

--Progress to next state
GenerateNextState:
process (CurrentState, DAV, CTS, full, empty)
	begin
		case CurrentState is
			when Start	=> if (DAV = '1' and full = '0') then
									NextState <= Write_memory;
								elsif (DAV = '0' and empty = '0' and CTS = '1') then
									NextState <= Attend_output;
								elsif (DAV = '1' and full = '1' and CTS = '1') then
									NextState <= Attend_output;
								else
									NextState <= Start;
								end if;
										
			when Write_memory	=> NextState <= Write_done;
									
								
			when Write_done => NextState <= IncrPut;
			
			
			when IncrPut => NextState <= Finish_write;
			
			
			when Finish_write => if (DAV = '0') then
											NextState <= Start;
										else
											NextState <= Finish_write;
										end if;
										
			when Attend_output => if (CTS = '0') then
											NextState <= Output_done;
										 else
											NextState <= Attend_output;
										 end if;
			
			when Output_done => NextState <= Start;
										 
		end case;
	end process;
	
--Output values
Wr <= '1' when(CurrentState = Write_done) else '0';
selnPG <= '1' when(CurrentState = Write_memory or CurrentState = Write_done or CurrentState = IncrPut) else '0';
incPut <= '1' when(CurrentState = IncrPut) else '0';
incGet <= '1' when(CurrentState = Output_done) else '0';
Wreg <= '1' when(CurrentState = Attend_output) else '0';
DAC <= '1' when(CurrentState = Finish_write) else '0';

end behavioral;